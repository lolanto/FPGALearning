`ifndef SIMPLE_CMD_EXECUTOR_V
`define SIMPLE_CMD_EXECUTOR_V

/**
 * 简易的命令执行器
 */

module SimpleCMDExecutor(
    input wire in_clk,
    input wire in_rst
);

endmodule

`endif // SMPLE_CMD_EXECUTOR_V