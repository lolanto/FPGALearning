module Top(
    input wire in_sig,
    output wire out_sig
);

    assign out_sig = in_sig;

endmodule
